-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Saturday, October 03, 2015 13:06:52 �й���׼ʱ��

